module changetoHex (
	input logic S0, S1, S2, S3, S4, S5, S6,
	output logic C0, C1, C2, C3, C4, C5, C6, C7, C8, C9, C10, C11
);


endmodule