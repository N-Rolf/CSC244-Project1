module changetoHex (
	input logic S0, S1, S2, S3, S4, S5, S6
	output logic C0, ... C11
);

	or (

endmodule