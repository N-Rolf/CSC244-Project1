module guffinOut_logic (
	input logic
	output logic
);



endmodule