module guffinOut_logic (
	input logic in_temp,
	output logic out_temp
);



endmodule